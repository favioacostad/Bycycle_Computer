`timescale 1ns / 1ps

module LCD_Bram_Big #(
    parameter RAM_WIDTH=8,
    parameter SYMBOL_WIDTH = 11,
    parameter LINEHEIGTH = 2
    )(
    input clock,
    input reset,
    input [14:0] address,
    input [2:0] enable,             //[0] = neuer Pixel-Schwung, [1] = neue Zeile, [2] = komplett neuer schreibprozess
    output [4:0] symbolwidth,
    output [RAM_WIDTH-1:0] out
    );
    
    reg [2:0] line;       
    assign symbolwidth = SYMBOL_WIDTH;
    reg [14:0]  address_ir;
    wire [10:0] address_iw;        
    assign address_iw = address_ir[10:0];
    reg [14:0] address_new;
    wire [14:0] ad;
    assign ad = ((1+address)*(LINEHEIGTH*SYMBOL_WIDTH))-1-(line*SYMBOL_WIDTH);       
    wire [7:0] data;    
    reg [7:0] data_int;    
    assign out = data_int;//address_ir > address_new - (SYMBOL_WIDTH)?data_int:8'd0;
    
    
    
    BRAM_SDP_MACRO #(
	    .BRAM_SIZE("18Kb"),             // Target BRAM, "18Kb" or "36Kb"
        .DEVICE("7SERIES"),             // Target device: "7SERIES"
        .WRITE_WIDTH(1),        // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(RAM_WIDTH),         // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .DO_REG(0),                     // Optional output register (0 or 1)
        .INIT_FILE("NONE"),
        .SIM_COLLISION_CHECK("ALL"),    // Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
        .SRVAL(72'd0),                  // Set/Reset value for port DO
        .INIT(72'd0),                   // Initial values on output port
        .WRITE_MODE("READ_FIRST"),      // Specify "READ_FIRST" for same clock or synchronous clocks, "WRITE_FIRST for asynchronous clocks on ports        
        .INIT_00(256'h0C101122222211100C0300000000000000000000000000000000000000000000),
        .INIT_01(256'hFECECFFFCFCEFEFCF0030F1F1E3D3D3D1E1F0F03F00C023231013132020CF003),
        .INIT_02(256'h03070F070301000000F0F8F8F0E0F0F8F8F00000000103070F0703010000F0FC),
        .INIT_03(256'hFCFCFCB8C0C080030707131B1F1B130707030080C0E0F0F8F0E0C08000000001),
        .INIT_04(256'h0000000000000080C0E0F0FCF0E0C08000000307171B1F1B1707030080C0C0B8),
        .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_07(256'h18780003070C08080C0703000000000000000000000000000000000000000000),
        .INIT_08(256'h0000000070F88C04048CF8700000000008093F3F0908000080C060202060C8A8),
        .INIT_09(256'h00060F0F07006078793F00000000000000000000000000000000000000000000),
        .INIT_0A(256'h80C8F030181E1830F0C880000907060C3C0C06070900000000FF3366CC98F000),
        .INIT_0B(256'h00000103070F1F0000000000FCF8F0E0C08000000000001F0F07030100000000),
        .INIT_0C(256'h10181CFE1C181000000000040C1C3F1C0C040000000080C0E0F0F8FC00000000),
        .INIT_0D(256'h00000000000000000000FEFE0000FEFE00000000003737000037370000000000),
        .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_1F(256'h0000000000383838000000000000000000000000000000000000000000000000),
        .INIT_20(256'h0000000080C0E070381C0E181C0E070301000000000000000000000000000000),
        .INIT_21(256'h003030303F3F30303000F8FE060383C363331EFEF8071F1E3331303030181F07),
        .INIT_22(256'h07030383C3E3773E1C30383C3E3733313030303000000C0C0EFFFF0000000000),
        .INIT_23(256'h030303033F3F03030C0E07C3C3C3C3C3E77E3C0C1C383030303030391F0E1C1E),
        .INIT_24(256'h63636363E3C3830C1C383030303030381F0FC0E070381C0E07FFFF0000030303),
        .INIT_25(256'h0F0300000000C0F0F8DCCEC7C3C3C380000F1F393030303030391F0F3F7F6363),
        .INIT_26(256'hC3E7FEBC000F1F393030303030391F0F030303030303C3F33F0F03000000303C),
        .INIT_27(256'h000000003C7EE7C3C3C3C3C3E7FEFC0000303030381C0E07030000BCFEE7C3C3),
        .INIT_28(256'h0000000000004E7E3E0000000000000000383838000000000000000007070700),
        .INIT_29(256'h0000000000000000000000000000000000000000000000000000003838380000),
        .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
               
        .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000) 
    ) BRAM_SDP_MACRO_inst (
        .DO(data), // Output read data port, width defined by READ_WIDTH parameter
        .DI(1'd0), // Input write data port, width defined by WRITE_WIDTH parameter
        .RDADDR(address_iw), // Input read address, width defined by read port depth
        .RDCLK(!clock), // 1-bit input read clock
        .RDEN(1'd1), // 1-bit input read port enable
        .REGCE(1'd0), // 1-bit input read output register enable
        .RST(reset), // 1-bit input reset
        .WE(1'd1), // Input write enable, width defined by write port depth
        .WRADDR(14'd0), // Input write address, width defined by write port depth
        .WRCLK(1'd0), // 1-bit input write clock
        .WREN(1'd0) // 1-bit input write port enable
    );
               
    always @(posedge clock) begin
        if(reset || enable[2]) begin
            address_new <= 0;
            address_ir  <= 0;
            data_int    <= 0;
            line        <= 0;
        end        
        else begin
            line <= line + enable[1];
            address_new <= ad; // address==0?address:ad;
            data_int <= address_ir > address_new-SYMBOL_WIDTH?data:8'd0;
            if(address_new != ad) begin             // if new address         
                address_ir <= ad;
            end
            else begin
                if(enable[0] && address_ir > address_new-SYMBOL_WIDTH)
                    address_ir <= address_ir - 1;
                else
                    address_ir <= address_ir;                    
            end
        end
    end      
    
endmodule
