`timescale 1ns / 1ps

module LCD_Bram_Small #(
    parameter RAM_WIDTH=8,
    parameter SYMBOL_WIDTH = 5,
    parameter LINEHEIGTH = 1
    )(
    input clock,
    input reset,
    input [14:0] address,
    input [2:0] enable,
    output [4:0] symbolwidth,
    output [RAM_WIDTH-1:0] out
    );
    
    
    reg [2:0] line;       
    assign symbolwidth = SYMBOL_WIDTH;
    reg [14:0]  address_ir;
    wire [10:0] address_iw;        
    assign address_iw = address_ir[10:0];


    reg [14:0] address_new;
    wire [14:0] ad;
    assign ad = ((1+address)*(LINEHEIGTH*SYMBOL_WIDTH))-1-(line*SYMBOL_WIDTH);    
    
    
    wire [7:0] data;    
    reg [7:0] data_int;    
    assign out = data_int;//address_ir > address_new - (SYMBOL_WIDTH)?data_int:8'd0;
    
    BRAM_SDP_MACRO #(
	    .BRAM_SIZE("18Kb"),             // Target BRAM, "18Kb" or "36Kb"
        .DEVICE("7SERIES"),             // Target device: "7SERIES"
        .WRITE_WIDTH(1),        // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(RAM_WIDTH),         // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .DO_REG(0),                     // Optional output register (0 or 1)
        .INIT_FILE("NONE"),
        .SIM_COLLISION_CHECK("ALL"),    // Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
        .SRVAL(72'd0),                  // Set/Reset value for port DO
        .INIT(72'd0),                   // Initial values on output port
        .WRITE_MODE("READ_FIRST"),      // Specify "READ_FIRST" for same clock or synchronous clocks, "WRITE_FIRST for asynchronous clocks on ports
      //.INIT_XX(256'h-->||<--05-->||<--04-->||<--03-->||<--02-->||<--01-->||<--00-->|),   
        .INIT_00(256'h5C1830367F3630183C7E3C181C3E7C3E1C3E6B6F6B3E3E4551453E0000000000),
      //.INIT_XX(256'h--0C-->||<--0B-->||<--0A-->||<--09-->||<--08-->||<--07-->||<--06), 
        .INIT_01(256'h2979290630484A360E0000000000000000000000000000000018180000185C7E),
        .INIT_02(256'h0014367F3614081C3E7F00007F3E1C082A1C361C2A607E0A353F000000000006),
        .INIT_03(256'h7F301004067F060414B6FFB6146060606000224D55592206097F017F005F005F),
        .INIT_04(256'h030F3F0F03303C3F3C30083E083E087840404040081C3E080808083E1C081030),
        .INIT_05(256'h20506313086463242B6A1200247E247E24070300070300065F06000000000000),
        .INIT_06(256'hE060000008083E0808083E1C3E0800413E0000003E4100000007030000364956),
        .INIT_07(256'h36625149494600427F40003E5149453E20100804020060600000080808080800),
        .INIT_08(256'h49291E364949493601710905033C4A4949302F494949311814127F1022494949),
        .INIT_09(256'h020159090600412214082424242424081422410000EC6C0000006C6C00000649),
        .INIT_0A(256'h09017F494949417F4141413E3E414141227F494949367E1111117E3E415D551E),
        .INIT_0B(256'h404040407F08142241304040403F00417F41007F0808087F3E4149497A7F0909),
        .INIT_0C(256'h327F090919663E4151215E7F090909063E4141413E7F0204087F7F0204027F7F),
        .INIT_0D(256'h70080763140814633F403C403F1F2040201F3F4040403F01017F010126494949),
        .INIT_0E(256'h808080808004020102040041417F000204081020007F41410071494543000708),
        .INIT_0F(256'h09003854545408384444447F38444444287F4444443820545454780003070000),
        .INIT_10(256'h007F40007F102844004080847D0000007D40007F0404780018A4A4A47C087E09),
        .INIT_11(256'h20447844040838444444FCFC4444443838444444387C040478007C0418047800),
        .INIT_12(256'h603C006C10106C003C6030603C1C2040201C3C40207C00043E44240008545454),
        .INIT_13(256'h003E4141413E0000007F0204087F0000007F0204027F0000007F404040400000),
        .INIT_14(256'h3C2623263C02010201000041413E080000770000083E4141006454544C009CA0),
        .INIT_15(256'h003F403C403F0000001F2040201F0000003F4040403F00000001017F01010000), /// <---------------
        .INIT_16(256'h00007F4141000000007149454300000000070870080700000063140814630000),
        .INIT_17(256'h80808080808000000004020102040000000041417F0000000002040810200000),
        .INIT_18(256'h0038444444280000007F44444438000000205454547800000000030700000000),
        .INIT_19(256'h0018A4A4A47C000000087E0909000000003854545408000000384444447F0000),
        .INIT_1A(256'h007F102844000000004080847D0000000000007D40000000007F040478000000),
        .INIT_1B(256'h0038444444380000007C040478000000007C0418047800000000007F40000000),
        .INIT_1C(256'h000854545420000000447844040800000038444444FC000000FC444444380000),
        .INIT_1D(256'h003C6030603C0000001C2040201C0000003C40207C00000000043E4424000000),
        .INIT_1E(256'h00083E4141000000006454544C000000009CA0603C000000006C10106C000000),
        .INIT_1F(256'h003C2623263C00000002010201000000000041413E0800000000007700000000),
        .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_21(256'h000000000000000000000000003333000000000000000000000000007CFFFF7C),
        .INIT_22(256'h000000000000000000000000000000003C000000000000000000003C3C00003C),
        .INIT_23(256'h030200000000000000021E1F03021E1FF07E1E100000000000001090F07E1E90),
        .INIT_24(256'h793F00000000000000060F0F0700307898F000000000000000000000FF3366CC),
        .INIT_25(256'h38383800000000000030381C0E070301E070381C0000000000003838380080C0),
        .INIT_26(256'h1C3622000000000000001F3F3121371E1C00000000000000000000B8FCC6E23E),
        .INIT_27(256'h00000000000000000000000000000000000000000000000000000000273F1F00),
        .INIT_28(256'h2000000000000000000000030F1F38200100000000000000000000F0FCFE0701),
        .INIT_29(256'h03000000000000000000002020381F0FF000000000000000000000010107FEFC),
        .INIT_2A(256'h0E0C00000000000000000C0E030F0F03B898000000000000000098B8E0F8F8E0),
        .INIT_2B(256'h010100000000000000000101010F0F0180800000000000000000808080F0F080),
        .INIT_2C(256'h000000000000000000000000B8F8780000000000000000000000000000000000),
        .INIT_2D(256'h0101000000000000000001010101010180800000000000000000808080808080),
        .INIT_2E(256'h0000000000000000000000003838380000000000000000000000000000000000),
        .INIT_2F(256'h000000000000000000181C0E0703010070381C0E00000000000000000080C0E0),
        .INIT_30(256'h30181F070000000000071F1E33313030331EFEF80000000000F8FE060383C363),
        .INIT_31(256'h30303000000000000000003030303F3F00000000000000000000000C0C0EFFFF),
        .INIT_32(256'h30303030000000000030383C3E373331E3773E1C00000000001C1E07030383C3),
        .INIT_33(256'h30391F0E00000000000C1C3830303030C3E77E3C00000000000C0E07C3C3C3C3),
        .INIT_34(256'h3F3F0303000000000003030303030303FFFF00000000000000C0E070381C0E07),
        .INIT_35(256'h30381F0F00000000000C1C383030303063E3C38300000000003F7F6363636363),
        .INIT_36(256'h30391F0F00000000000F1F3930303030C3C380000000000000C0F0F8DCCEC7C3),
        .INIT_37(256'h000000000000000000000000303C0F03F33F0F030000000000030303030303C3),
        .INIT_38(256'h30391F0F00000000000F1F3930303030E7FEBC00000000000000BCFEE7C3C3C3),
        .INIT_39(256'h0E07030000000000000000303030381CC3E7FEFC00000000003C7EE7C3C3C3C3),
        .INIT_3A(256'h0000000000000000000000001C1C1C0000000000000000000000000070707000),
        .INIT_3B(256'h0000000000000000000000009CFC7C0000000000000000000000000070707000),
        .INIT_3C(256'h38300000000000000000000103070E1C07030000000000000000C0E0F0381C0E),
        .INIT_3D(256'h0606060000000000000006060606060660606000000000000000606060606060),
        .INIT_3E(256'h0100000000000000000030381C0E0703E0C0000000000000000003070E1C38F0),
        .INIT_3F(256'h00000000000000000000000000373700773E1C0000000000001C1E070383C3E3),
        // The next set of INIT_xx are valid when configured as 36Kb
        .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000) 
    ) BRAM_SDP_MACRO_inst (
        .DO(data), // Output read data port, width defined by READ_WIDTH parameter
        .DI(1'd0), // Input write data port, width defined by WRITE_WIDTH parameter
        .RDADDR(address_iw), // Input read address, width defined by read port depth
        .RDCLK(!clock), // 1-bit input read clock
        .RDEN(1'd1), // 1-bit input read port enable
        .REGCE(1'd0), // 1-bit input read output register enable
        .RST(reset), // 1-bit input reset
        .WE(1'd1), // Input write enable, width defined by write port depth
        .WRADDR(14'd0), // Input write address, width defined by write port depth
        .WRCLK(1'd0), // 1-bit input write clock
        .WREN(1'd0) // 1-bit input write port enable
    );
     
    always @(posedge clock) begin
       if(reset || enable[2]) begin
           address_new <= 0;
           address_ir  <= 0;
           data_int    <= 0;
           line        <= 0;
       end        
       else begin
           line <= line + enable[1];
           address_new <= ad; // address==0?address:ad;
           data_int <= address_ir > address_new-SYMBOL_WIDTH?data:8'd0;
           if(address_new != ad) begin             // if new address         
               address_ir <= ad;
           end
           else begin
               if(enable[0] && address_ir > address_new-SYMBOL_WIDTH)
                   address_ir <= address_ir - 1;
               else
                   address_ir <= address_ir;                    
           end
       end
    end 
        
    /*   
    always @(posedge clock) begin
        if(reset) begin
            address_new <= 0;
            address_ir  <= 0;
            data_int    <= 0;
        end        
        else begin
            address_new <= ad; // address==0?address:ad;
            data_int <= address_ir > address_new-SYMBOL_WIDTH?data:8'd0;
            if(address_new != ad) begin             // if new address         
                address_ir <= ad;
            end
            else begin
                if(enable[0] && address_ir > address_new-SYMBOL_WIDTH)
                    address_ir <= address_ir - 1;
                else
                    address_ir <= address_ir;                    
            end
        end
    end    
    */
endmodule
